library verilog;
use verilog.vl_types.all;
entity tbDatapath is
end tbDatapath;

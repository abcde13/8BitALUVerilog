library verilog;
use verilog.vl_types.all;
entity tbMain is
end tbMain;

library verilog;
use verilog.vl_types.all;
entity tbControl is
end tbControl;

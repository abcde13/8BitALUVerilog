library verilog;
use verilog.vl_types.all;
entity subtractor is
    port(
        cin             : in     vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic;
        cout            : out    vl_logic;
        z               : out    vl_logic
    );
end subtractor;
